// =============================================================================
//  rk4_uart_sequencer.sv -- UVM sequencer for UART TX items
// =============================================================================
typedef uvm_sequencer #(rk4_uart_tx_item) rk4_uart_sequencer;
